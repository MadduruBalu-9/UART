`include "uvm_macros.svh"
 import uvm_pkg::*;


`include "uart_if.sv"
`include "uart_seq_item.sv"

//Sequences
`include "rand_baud.sv"

//Driver

`include "driver.sv"

//Monitor

//`include "mon.sv"

//Agent.sv

`include "agent.sv"


//Sco

//`include "sco.sv"

//Env

`include "env.sv"

//test

`include "test.sv"

